library verilog;
use verilog.vl_types.all;
entity div_32bit_tb is
end div_32bit_tb;

`timescale 1ns/ 1ps

module multiplexer32to1_tb;
    
    // Inputs
    reg [31:0] BusMuxIn_R0;
    reg [31:0] BusMuxIn_R1;
    reg [31:0] BusMuxIn_R2;
    reg [31:0] BusMuxIn_R3; 
    reg [31:0] BusMuxIn_R4;
    reg [31:0] BusMuxIn_R5;
    reg [31:0] BusMuxIn_R6;
    reg [31:0] BusMuxIn_R7;
    reg [31:0] BusMuxIn_R8;
    reg [31:0] BusMuxIn_R9;
    reg [31:0] BusMuxIn_R10;
    reg [31:0] BusMuxIn_R11;
    reg [31:0] BusMuxIn_R12;
    reg [31:0] BusMuxIn_R13;
    reg [31:0] BusMuxIn_R14;
    reg [31:0] BusMuxIn_R15;
    reg [31:0] BusMuxIn_HI;
    reg [31:0] BusMuxIn_LO;
    reg [31:0] BusMuxIn_Z_high;
    reg [31:0] BusMuxIn_Z_low;
    reg [31:0] BusMuxIn_PC;
    reg [31:0] BusMuxIn_MDR;    
    reg [31:0] BusMuxIn_InPort;
    reg [31:0] C_sign_extended;
    reg [31:0] BusMuxIn_Y;
    reg [4:0] select_signal;
    
    // Output
    wire [31:0] BusMuxOut;

endmodule
library verilog;
use verilog.vl_types.all;
entity mul_32bit_tb is
end mul_32bit_tb;

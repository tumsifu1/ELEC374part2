library verilog;
use verilog.vl_types.all;
entity storeTB is
end storeTB;

library verilog;
use verilog.vl_types.all;
entity sub_32tb is
end sub_32tb;

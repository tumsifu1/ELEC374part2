library verilog;
use verilog.vl_types.all;
entity shr_TB is
end shr_TB;

library verilog;
use verilog.vl_types.all;
entity bidirectional_bus is
    port(
        R0Signal        : in     vl_logic;
        R1Signal        : in     vl_logic;
        R2Signal        : in     vl_logic;
        R3Signal        : in     vl_logic;
        R4Signal        : in     vl_logic;
        R5Signal        : in     vl_logic;
        R6Signal        : in     vl_logic;
        R7Signal        : in     vl_logic;
        R8Signal        : in     vl_logic;
        R9Signal        : in     vl_logic;
        R10Signal       : in     vl_logic;
        R11Signal       : in     vl_logic;
        R12Signal       : in     vl_logic;
        R13Signal       : in     vl_logic;
        R14Signal       : in     vl_logic;
        R15Signal       : in     vl_logic;
        HISignal        : in     vl_logic;
        LOSignal        : in     vl_logic;
        ZHISignal       : in     vl_logic;
        ZLOSignal       : in     vl_logic;
        PCSignal        : in     vl_logic;
        MDRSignal       : in     vl_logic;
        InportSignal    : in     vl_logic;
        CSignal         : in     vl_logic;
        encoderY        : in     vl_logic;
        BusMuxInputs_R0 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R1 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R2 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R3 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R4 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R5 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R6 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R7 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R8 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R9 : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R10: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R11: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R12: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R13: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R14: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_R15: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_HI : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_LO : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_Z_high: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_Z_low: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_PC : in     vl_logic_vector(31 downto 0);
        BusMuxInputs_MDR: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_InPort: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_C_sign_extended: in     vl_logic_vector(31 downto 0);
        BusMuxInputs_Y  : in     vl_logic_vector(31 downto 0);
        BusMuxOutToDatapath: out    vl_logic_vector(31 downto 0)
    );
end bidirectional_bus;

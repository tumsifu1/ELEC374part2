library verilog;
use verilog.vl_types.all;
entity MDRTB is
end MDRTB;

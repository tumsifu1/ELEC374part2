library verilog;
use verilog.vl_types.all;
entity div_tb is
end div_tb;

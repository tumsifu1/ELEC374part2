library verilog;
use verilog.vl_types.all;
entity add_TB is
end add_TB;
